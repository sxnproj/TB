interface if_dft;

    var logic scan_en;
    var logic test_mode;
    var logic scan_in0;
    var logic scan_out0;

endinterface : if_dft