package usbf_top_pkg;
    import uvm_pkg::*;

    `include "src/uvm/sequence_items/packet_transaction.sv"
    `include "src/uvm/sequence_items/packet_init.sv"
    `include "src/uvm/sequence_items/endpoint_data.sv"
    `include "src/uvm/sequence_items/interrupt_data.sv"
    `include "src/uvm/sequence_items/func_address.sv"
    `include "src/uvm/sequence_items/buffer_size.sv"
    `include "src/uvm/sequence_items/packet_data.sv"
    `include "src/uvm/sequence_items/wb_read_data.sv"
    `include "src/uvm/sequence_items/utmi_read_data.sv"
    `include "src/uvm/sequence_transaction.sv"
    `include "src/uvm/subscribers/endpoint_data_sub.sv"
    `include "src/uvm/subscribers/packet_init_sub.sv"
    `include "src/uvm/subscribers/packet_transaction_sub.sv"
    `include "src/uvm/subscribers/interrupt_data_sub.sv"
    `include "src/uvm/subscribers/func_address_sub.sv"
    `include "src/uvm/subscribers/buffer_size_sub.sv"
    `include "src/uvm/subscribers/packet_data_sub.sv"
    `include "src/uvm/subscribers/wb_done_sub.sv"
    `include "src/uvm/subscribers/utmi_done_sub.sv"
    `include "src/uvm/subscribers/data_buffer_sub.sv"
    `include "src/uvm/subscribers/wb_data_sub.sv"
    `include "src/uvm/subscribers/utmi_data_sub.sv"
    `include "src/uvm/sequence_init.sv"
    `include "src/uvm/sequencer_transaction.sv"
    `include "src/uvm/sequencer_init.sv"
    `include "src/uvm/sequencer_virtual.sv"
    `include "src/uvm/sequence_virtual.sv"
    `include "src/uvm/driver_utmi.sv"
    `include "src/uvm/driver_wb.sv"
    `include "src/uvm/monitor_utmi.sv"
    `include "src/uvm/monitor_wb.sv"
    `include "src/uvm/agent_utmi.sv"
    `include "src/uvm/agent_wb.sv"
    `include "src/uvm/env.sv"
    `include "src/usbf_top_test.sv"

endpackage : usbf_top_pkg